// BMP280.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module BMP280 (
		output wire [31:0] address,       // avalon_master.address
		output wire        read,          //              .read
		input  wire [31:0] readdata,      //              .readdata
		input  wire        readdatavalid, //              .readdatavalid
		input  wire        waitrequest,   //              .waitrequest
		output wire        write,         //              .write
		output wire [3:0]  byteenable,    //              .byteenable
		output wire [31:0] writedata,     //              .writedata
		input  wire        clk,           //         clock.clk
		input  wire        i2c_data_in,   //   conduit_end.conduit_data_in
		input  wire        i2c_clk_in,    //              .conduit_clk_in
		output wire        i2c_data_oe,   //              .conduit_data_oe
		output wire        i2c_clk_oe,    //              .conduit_clk_oe
		input  wire        rst_n          //         reset.reset_n
	);

	altera_i2cslave_to_avlmm_bridge #(
		.I2C_SLAVE_ADDRESS (7'b1110111),
		.BYTE_ADDRESSING   (1),
		.ADDRESS_STEALING  (0),
		.READ_ONLY         (0)
	) i2cslave_to_avlmm_bridge_0 (
		.clk           (clk),           //         clock.clk
		.address       (address),       // avalon_master.address
		.read          (read),          //              .read
		.readdata      (readdata),      //              .readdata
		.readdatavalid (readdatavalid), //              .readdatavalid
		.waitrequest   (waitrequest),   //              .waitrequest
		.write         (write),         //              .write
		.byteenable    (byteenable),    //              .byteenable
		.writedata     (writedata),     //              .writedata
		.rst_n         (rst_n),         //         reset.reset_n
		.i2c_data_in   (i2c_data_in),   //   conduit_end.conduit_data_in
		.i2c_clk_in    (i2c_clk_in),    //              .conduit_clk_in
		.i2c_data_oe   (i2c_data_oe),   //              .conduit_data_oe
		.i2c_clk_oe    (i2c_clk_oe)     //              .conduit_clk_oe
	);

endmodule
